----------------------------------------------------------------------------------
-- Company: 
-- Engineer: Javier Antonio Ricaldi Esquivel
--           Dario Fernando Gallegos Quispe
-- 
-- Create Date:    15:08:40 05/25/2018 
-- Design Name: 
-- Module Name:    ram2 - syn 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity ram2 is
  port ( 
    rst_n : in  std_logic;   -- reset asíncrono del sistema (a baja)
    clk   : in  std_logic;   -- reloj del sistema
	 dInB 	: in  std_logic_vector (3 downto 0);
	 addrA	: in  std_logic_vector (14 downto 0);
	 addrB : in std_logic_vector (14 downto 0);
	 weB	: in  std_logic;
	 dOutA 	: out std_logic_vector (3 downto 0);
	 dOutB 	: out std_logic_vector (3 downto 0)
    );
end ram2;

use work.common.all;

architecture syn of ram2 is

	constant	DATA_WIDTH	: natural := 4;
	constant MAX_SIZE		: natural := 19_200;

	type ramType is array (0 to MAX_SIZE -1) of std_logic_vector (DATA_WIDTH - 1 downto 0);
  signal ram : ramType := (X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"7",X"7",X"7",X"7",X"7",X"7",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",X"4",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"B",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"f",X"7",X"7",X"7",X"7",X"7",X"7",X"f",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",X"8",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",
									X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7",X"7");
  


begin

	lecturaCampo:
	process (clk)
	begin
		if rising_edge(clk) then
				dOutA <= ram( to_integer( unsigned( addrA ) ) ) ;
		end if;
	end process;
	
	rw:
	process (clk)
	begin
		if rising_edge(clk) then
			if weB='1' then
				ram(to_integer(unsigned( addrB ) ) ) <= dInB;
			else
				dOutB <= ram( to_integer( unsigned( addrB ) ) ) ;
				
			end if;
		end if;
	end process;

end syn;

